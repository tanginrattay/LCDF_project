// File: top.sv
// Description: Top-level module for the game. Connects all sub-modules for
//              game logic, map generation, and VGA output.
// --- THIS FILE CONTAINS THE CRITICAL FIX ---

module top(
    input wire clk,         // Main input clock (e.g., 100MHz)
    input wire RST_n,       // On-board reset button (active-low)
    input wire [2:0] sw,    // Switches for game control
    output wire [3:0] R,    // VGA Red output
    output wire [3:0] G,    // VGA Green output
    output wire [3:0] B,    // VGA Blue output
    output wire HS,         // VGA Horizontal Sync
    output wire VS,         // VGA Vertical Sync
//    output wire beep,
    output wire [1:0] gamemode_led
);

    // --- Internal Signals ---
    wire rst_n_debounced; // Debounced active-low reset signal
    wire clk_25mhz;       // 25MHz clock for VGA pixel timing
    wire clk_60hz;        // 60Hz clock for game logic timing
    
    wire [1:0] gamemode;
    wire [8:0] player_y;

    // SystemVerilog arrays (busses) to connect modules
    logic [9:0] [19:0] obstacle_x_bus;
    logic [9:0] [17:0] obstacle_y_bus;

    // VGA signals
    wire [9:0] pix_x;
    wire [8:0] pix_y;
    wire [11:0] vga_data_out; // 12-bit color data from screen generator

    // --- Debouncer Instantiation ---
    // *** CRITICAL FIX: This was missing. ***
    // This module creates a clean, debounced reset signal from the physical button.
    // Assuming your module is named Anti_jitter. If not, replace the name.
    // Anti_jitter u_anti_jitter (.clk(clk), .rst_in(RST_n), .rst_out(rst_n_debounced));
    // If you don't have a debouncer, for now, you can bypass it to test:
    assign rst_n_debounced = RST_n;


    // --- Clock Generation ---
    // Generate 25MHz clock for VGA from main clock (assuming 100MHz input)
    reg [1:0] clk_div_25m;
    always_ff @(posedge clk or negedge rst_n_debounced) begin
        if (!rst_n_debounced) clk_div_25m <= 2'b0;
        else clk_div_25m <= clk_div_25m + 1;
    end
    assign clk_25mhz = clk_div_25m[1];

    // Generate 60Hz clock for game logic
    // Assuming you have a module named clkdiv_60hz
    clkdiv_60hz u_clkdiv_60hz(.clk(clk), .rst_n(rst_n_debounced), .clk_60hz(clk_60hz));


    // --- Game Logic Module ---
    game_logic u_game_logic (
        .rst_n(rst_n_debounced),
        .sw(sw),
        .clk(clk_60hz),
        .obstacle_x(obstacle_x_bus),
        .obstacle_y(obstacle_y_bus),
        .gamemode(gamemode),
        .player_y(player_y)
    );

    // --- Map Generation Module ---
    map u_map (
        .rst_n(rst_n_debounced),
        .clk(clk_60hz),
        .gamemode(gamemode),
        .obstacle_x(obstacle_x_bus),
        .obstacle_y(obstacle_y_bus)
    );

    // --- VGA Screen Picture Generator ---
    vga_screen_pic u_vga_screen_pic(
        .pix_x(pix_x),
        .pix_y(pix_y),
        .gamemode(gamemode),
        .player_y(player_y),
        .obstacle_x(obstacle_x_bus),
        .obstacle_y(obstacle_y_bus),
        .rgb(vga_data_out)
    );

    // --- VGA Controller ---
    // This module generates the HS/VS sync signals and outputs the final color data.
    // Assuming you have a module named vga_ctrl
    vga_ctrl u_vga_ctrl(
        .clk(clk_25mhz),
        .rst(~rst_n_debounced), // vga_ctrl often uses an active-high reset
        .Din(vga_data_out),
        .row(pix_y),
        .col(pix_x),
        // .rdn(rdn), // This signal is generated by vga_ctrl but not used elsewhere
        .R(R),
        .G(G),
        .B(B),
        .HS(HS),
        .VS(VS)
    );
    
    // --- Other Peripherals ---
    assign gamemode_led = gamemode;

    // Assuming you have a module named top_beep
//    top_beep u_top_beep(
//        .clk(clk),
//        .gamemode(gamemode),
//        .beep(beep)
//    );

endmodule